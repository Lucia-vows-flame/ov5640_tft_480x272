module ov5640_tft_480x272
(
        input                   i_sysclk                , // system clock
        input                   i_sysrst_n              , // system reset
        // camera interface
        input                   i_ov5640_pclk           , // camera pixel clock
        input                   i_ov5640_vsync          , // camera vsync signal
        input                   i_ov5640_href           , // camera href signal
        input       [7:0]       i_ov5640_data           , // camera data
        output                  camera_rst_n            , // camera reset signal
        output                  camera_pwdn             , // camera power down signal
        output                  sccb_scl                , // sccb clock signal
        inout                   sccb_sda                , // sccb data signal
        // sdram interface
        output                  sdram_clk               , // sdram clock
        output                  sdram_cke               , // sdram clock enable
        output                  sdram_cs_n              , // sdram chip select
        output                  sdram_ras_n             , // sdram row address select
        output                  sdram_cas_n             , // sdram column address select
        output                  sdram_we_n              , // sdram write enable
        output      [1:0]       sdram_ba                , // sdram bank address
        output      [12:0]      sdram_addr              , // sdram address
        inout       [15:0]      sdram_dq                , // sdram data
        output      [1:0]       sdram_dqm               , // sdram data mask
        // tft interface
        output                  o_tft_clk               , // tft pixel clock
        output                  o_tft_de                , // tft data enable
        output                  o_tft_bl                , // tft backlight control
        output                  o_tft_hsync             , // tft hsync signal
        output                  o_tft_vsync             , // tft vsync signal
        output      [15:0]      o_tft_rgb_data            // tft rgb data
);

//********************************Parameter********************************//
parameter       H_PIXEL = 24'd480       ; // tft pixel width, used to set sdram cache size
parameter       V_PIXEL = 24'd272       ; // tft pixel height, used to set sdram cache size

//********************************Internal Wire and Reg define**************************//
// wire define
wire            clk_100m                ; // 100 MHz clock
wire            clk_100m_shift          ; // 100 MHz clock with phase shift
wire            clk_9m                  ; // 9 MHz clock
wire            sys_rst_n               ; // system reset
wire            camera_init_done        ; // camera init done signal
wire            wr_req                  ; // sdram write request
wire    [15:0]  wr_data                 ; // sdram write data
wire            rd_req                  ; // sdram read request, rd_req is generated by tft_disp module
wire    [15:0]  rd_data                 ; // sdram read data
wire            sdram_init_done         ; // sdram init done signal
wire            sys_init_done           ; // system init done signal : camera init done and sdram init done

//*****************************Main Code************************************//
// sys_init_done
assign  sys_init_done = camera_init_done & sdram_init_done;

//****************************Instantiation****************************//
// clk_and_rst
clk_and_rst u_clk_and_rst(
        .i_clk      	(i_sysclk       ),
        .i_rst_n    	(i_sysrst_n     ),
        .clk_9m     	(clk_9m         ),
        .clk_100m   	(clk_100m       ),
        .clk_100m_2 	(clk_100m_shift ),
        .sys_rst_n  	(sys_rst_n      )
);

// ov5640_top
ov5640_top u_ov5640_top(
        .i_sysclk         	(clk_9m            ),
        .i_pclk           	(i_ov5640_pclk     ),
        .i_sysrst_n       	(sys_rst_n         ),
        .i_vsync          	(i_ov5640_vsync    ),
        .i_href           	(i_ov5640_href     ),
        .i_data           	(i_ov5640_data     ),
        .i_sys_init_done  	(sys_init_done     ),
        .data_valid       	(wr_req            ), // data valid signal is used to control sdram fifo write enable
        .rgb_data         	(wr_data           ),
        .camera_init_done 	(camera_init_done  ),
        .camera_rst_n     	(camera_rst_n      ),
        .camera_pwdn      	(camera_pwdn       ),
        .iic_sclk         	(sccb_scl          ),
        .iic_sdat         	(sccb_sda          )
);

// sdram_top
sdram_top u_sdram_top(
        // system port
        .i_sysclk        	(clk_100m         ),
        .sdram_clk_in    	(clk_100m_shift   ),
        .i_sysrst_n      	(sys_rst_n        ),
        // user write port
        .wr_fifo_wr_clk  	(i_ov5640_pclk    ), // ov5640 writes data to fifo, so fifo write clock is ov5640 pclk
        .wr_fifo_wr_req  	(wr_req           ), // ov5640 data valid signal is used to control sdram fifo write enable
        .wr_fifo_wr_data 	(wr_data          ), // ov5640 data output is used for sdram write data
        .sdram_wr_b_addr 	(24'd0            ), // sdram write start address is 0
        .sdram_wr_e_addr 	(H_PIXEL * V_PIXEL), // sdram write end address is H_PIXEL * V_PIXEL
        .wr_burst_len    	(10'd512          ), // sdram burst length is 512
        .wr_rst          	(!sys_rst_n       ), // sys_rst_n is used to reset sdram fifo, but note that the reset signal of fifo is high level valid
        // user read port
        .rd_fifo_rd_clk  	(clk_9m           ), // tft read data from fifo, so fifo read clock is tft clk
        .rd_fifo_rd_req  	(rd_req           ), // rd_req is generated by tft_disp module
        .sdram_rd_b_addr 	(24'd0            ), // sdram read start address is 0
        .sdram_rd_e_addr 	(H_PIXEL * V_PIXEL), // sdram read end address is H_PIXEL * V_PIXEL
        .rd_burst_len    	(10'd512          ), // sdram burst length is 512
        .rd_rst          	(!sys_rst_n       ), // sys_rst_n is used to reset sdram fifo, but note that the reset signal of fifo is high level valid
        .rd_fifo_rd_data 	(rd_data          ), // sdram read data output
        .rd_fifo_num     	(                 ), // In this design, rd_fifo_num is not used, so it is not connected
        // user control port
        .read_valid      	(1'b1             ), // read valid signal is always high
        .init_end        	(sdram_init_done  ), // sdram init done signal
        .pingpang_enable 	(1'b1             ), // pingpang enable signal is always high, because we use pingpang mode
        .sdram_clk_out   	(sdram_clk        ),
        .sdram_cke       	(sdram_cke        ),
        .sdram_cs_n      	(sdram_cs_n       ),
        .sdram_ras_n     	(sdram_ras_n      ),
        .sdram_cas_n     	(sdram_cas_n      ),
        .sdram_we_n      	(sdram_we_n       ),
        .sdram_ba        	(sdram_ba         ),
        .sdram_addr      	(sdram_addr       ),
        .sdram_dqm       	(sdram_dqm        ),
        .sdram_dq        	(sdram_dq         )
);

// tft_disp
tft_disp u_tft_disp(
        .i_clk_9m      	(clk_9m         ),
        .i_sysrst_n    	(sys_rst_n      ),
        .i_data_in     	(rd_data        ), // The data of tft_disp comes from the data read out by read fifo
        .read_data_req 	(read_req       ), // read_req is generated by tft_disp module
        .rgb_data_tft  	(o_tft_rgb_data ), // tft rgb data output
        .tft_hsync     	(o_tft_hsync    ),
        .tft_vsync     	(o_tft_vsync    ),
        .tft_clk       	(o_tft_clk      ),
        .tft_de        	(o_tft_de       ),
        .tft_bl        	(o_tft_bl       )
);

endmodule